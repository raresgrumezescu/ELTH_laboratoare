R1	0 1 2
R2	3 1 1
R3	1 2 4
R5	3 4 2
H2 2 1 V1 2
V1	4 0 12	
V3	2 3 4
J4	1 4 4
*
.OP
.PRINT DC I(R1) I(R2) I(R3) I(R5) V(J4)
.END

