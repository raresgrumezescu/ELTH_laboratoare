R1 2 1 2
R2 4 3 2
R3 2 4 2
R4 4 5 2
V1 1 5 12
V2 3 2 6
G5 4 5 2 1 1
.OP
.PRINT DC I(R1) I(R2) I(R3) I(R4) I(G5)
.END
