*
R1 1 2 5
R3 2 3 4
R4 4 5 3
R5 5 4 2
V1 5 1 78
E3 3 5 5 2 0.5
F5 5 2 V4 0.5
V4 2 6 0
*
.OP
.PRINT DC I(R1) I(R3) I(R4) I(R5) I(F5)
.END
